module imm_gen.sv ();
endmodule