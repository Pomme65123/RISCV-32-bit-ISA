module instr_memory.sv ();
endmodule