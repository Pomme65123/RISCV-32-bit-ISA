module hazard_detection_unit ();
endmodule