module alu ();
endmodule