module riscv_cpu_tb ();
endmodule